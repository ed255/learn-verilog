// Binary add
module main (
  input wire [5:0] a,
  input wire [5:0] b,
  output wire [5:0] c
);

  assign c = a / b;

endmodule

